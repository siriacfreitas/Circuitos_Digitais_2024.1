LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY Lab_04_linha3 is 
    PORT(
         NUM3: in std_logic_vector(3 downto 0);
         LINHA3: out std_logic_vector (7 downto 0);
        );
END ENTITY;

ARCHITECTURE main OF Lab_04_linha3 is
    begin
        LINHA3(0) <= '0'
        LINHA3(1) <= (NOT(NUM3(2)) AND NOT(NUM3(1)) AND NOT(NUM3(0))) OR (NOT(NUM3(2) AND NUM3(1) AND NUM3(0))) OR (NUM3(2) AND NOT(NUM3(1)) AND NUM3(0)) OR (NOT(NUM3(3)) AND NUM3(2) AND NOT(NUM3(0))) OR (NOT(NUM3(1)) AND NUM3(3));
        LINHA3(2) <= (NOT(NUM3(3)) AND NUM3(2) AND NOT(NUM3(1)) AND NOT(NUM3(0))) OR  (NUM3(3) AND NOT(NUM3(2)) AND NUM3(1) AND NOT(NUM3(0)));
        LINHA3(3) <= (NOT(NUM3(3)) AND NOT(NUM3(2)) AND NOT(NUM3(1)) AND NUM3(0)) OR  (NUM3(3) AND NUM3(2) AND NUM3(1) AND NUM3(0));
        LINHA3(4) <= (NOT(NUM3(3)) AND NUM3(2) AND NUM3(1) AND NUM3(0));
        LINHA3(5) <= (NOT(NUM3(2)) AND NOT(NUM3(0))) OR (NOT(NUM3(2)) AND NUM3(1)) OR (NUM3(1) AND NOT(NUM(0))) OR (NUM3(2) AND NOT(NUM3(1)) AND NUM3(0)) OR (NUM3(3) AND NOT(NUM3(0)));
        LINHA3(6) <= '0';
        LINHA3(7) <= '0';

END ARCHITECTURE;





LINHA6(0) <= 0

LINHA6(1) <= (NOT (NUM(3)) AND NUM6(2) AND NUM6(0)) OR (NUM6(2) AND NOT NUM6(1) AND NUM6(0))

LINHA6(2) <= (NOT (NUM6(3)) AND NOT (NUM6(0))) OR (NOT (NUM6(3)) AND NUM6(1)) OR (NOT (NUM6(3)) AND NUM6(2)) OR (NUM6(2) AND  NUM6(1) AND  NUM6(0)) OR (NUM6(3)) AND  NOT (NUM6(2)) AND NOT (NUM6(1))

LINHA6(3) <= (NOT (NUM6(2)) AND NOT (NUM6(1)) OR (NOT (NUM6(3)) AND NUM60) OR (NOT (NUM6(3))  AND NUM6(1))

LINHA6(4) <= (NOT (NUM6(3)) AND NOT (NUM6(2)) AND  NOT (NUM6(0))) OR (NOT (NUM6(3)) AND  NOT (NUM6(2)) AND  NUM6(1))) OR  (NOT (NUM6(3)) AND  NUM6(2) AND  NUM6(0)) OR (NUM6(3)  AND NOT (NUM6(2)) AND  NOT (NUM6(1)))

LINHA6(5) <=  (NOT (NUM6(3)) AND  NUM6(2) AND  NUM6(0)) OR (NUM6(3) AND  NOT (NUM6(2)) AND  NUM6(1) AND  NUM6(0))

LINHA3(6) <= '0';
LINHA3(7) <= '0';